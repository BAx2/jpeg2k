// Created with Corsair v1.0.2.dev0+894dec23

`ifndef __DMAREGS_VH
`define __DMAREGS_VH

`define DMA_CSR_BASE_ADDR 0
`define DMA_CSR_DATA_WIDTH 32
`define DMA_CSR_ADDR_WIDTH 8

// DEBUG_CR - DMA Control
`define DMA_CSR_DEBUG_CR_ADDR 8'hf0
`define DMA_CSR_DEBUG_CR_RESET 32'h0

// DEBUG_CR.MM2S_LEN - The burst length
`define DMA_CSR_DEBUG_CR_MM2S_LEN_WIDTH 8
`define DMA_CSR_DEBUG_CR_MM2S_LEN_LSB 0
`define DMA_CSR_DEBUG_CR_MM2S_LEN_MASK 32'hf0
`define DMA_CSR_DEBUG_CR_MM2S_LEN_RESET 8'h0

// DEBUG_CR.MM2S_SIZE - The number of bytes in a transfer must be equal to the data bus width
`define DMA_CSR_DEBUG_CR_MM2S_SIZE_WIDTH 3
`define DMA_CSR_DEBUG_CR_MM2S_SIZE_LSB 8
`define DMA_CSR_DEBUG_CR_MM2S_SIZE_MASK 32'hf0
`define DMA_CSR_DEBUG_CR_MM2S_SIZE_RESET 3'h0

// DEBUG_CR.MM2S_START - Start read transaction
`define DMA_CSR_DEBUG_CR_MM2S_START_WIDTH 1
`define DMA_CSR_DEBUG_CR_MM2S_START_LSB 12
`define DMA_CSR_DEBUG_CR_MM2S_START_MASK 32'hf0
`define DMA_CSR_DEBUG_CR_MM2S_START_RESET 1'h0

// DEBUG_CR.S2MM_LEN - The burst length
`define DMA_CSR_DEBUG_CR_S2MM_LEN_WIDTH 8
`define DMA_CSR_DEBUG_CR_S2MM_LEN_LSB 16
`define DMA_CSR_DEBUG_CR_S2MM_LEN_MASK 32'hf0
`define DMA_CSR_DEBUG_CR_S2MM_LEN_RESET 8'h0

// DEBUG_CR.S2MM_SIZE - The number of bytes in a transfer must be equal to the data bus width
`define DMA_CSR_DEBUG_CR_S2MM_SIZE_WIDTH 3
`define DMA_CSR_DEBUG_CR_S2MM_SIZE_LSB 24
`define DMA_CSR_DEBUG_CR_S2MM_SIZE_MASK 32'hf0
`define DMA_CSR_DEBUG_CR_S2MM_SIZE_RESET 3'h0

// DEBUG_CR.S2MM_START - Start read transaction
`define DMA_CSR_DEBUG_CR_S2MM_START_WIDTH 1
`define DMA_CSR_DEBUG_CR_S2MM_START_LSB 28
`define DMA_CSR_DEBUG_CR_S2MM_START_MASK 32'hf0
`define DMA_CSR_DEBUG_CR_S2MM_START_RESET 1'h0


// DEBUG_SR - DMA Status
`define DMA_CSR_DEBUG_SR_ADDR 8'hf4
`define DMA_CSR_DEBUG_SR_RESET 32'h0

// DEBUG_SR.MM2S_BUSY - Read transaction in process
`define DMA_CSR_DEBUG_SR_MM2S_BUSY_WIDTH 1
`define DMA_CSR_DEBUG_SR_MM2S_BUSY_LSB 0
`define DMA_CSR_DEBUG_SR_MM2S_BUSY_MASK 32'hf4
`define DMA_CSR_DEBUG_SR_MM2S_BUSY_RESET 1'h0

// DEBUG_SR.S2MM_BUSY - Write transaction in process
`define DMA_CSR_DEBUG_SR_S2MM_BUSY_WIDTH 1
`define DMA_CSR_DEBUG_SR_S2MM_BUSY_LSB 1
`define DMA_CSR_DEBUG_SR_S2MM_BUSY_MASK 32'hf4
`define DMA_CSR_DEBUG_SR_S2MM_BUSY_RESET 1'h0


// DEBUG_MM2S_ADDR - MM2S Start address
`define DMA_CSR_DEBUG_MM2S_ADDR_ADDR 8'hf8
`define DMA_CSR_DEBUG_MM2S_ADDR_RESET 32'h0

// DEBUG_MM2S_ADDR.ADDR - Indicates the Start Address
`define DMA_CSR_DEBUG_MM2S_ADDR_ADDR_WIDTH 32
`define DMA_CSR_DEBUG_MM2S_ADDR_ADDR_LSB 0
`define DMA_CSR_DEBUG_MM2S_ADDR_ADDR_MASK 32'hf8
`define DMA_CSR_DEBUG_MM2S_ADDR_ADDR_RESET 32'h0


// DEBUG_S2MM_ADDR - S2MM Start address
`define DMA_CSR_DEBUG_S2MM_ADDR_ADDR 8'hfc
`define DMA_CSR_DEBUG_S2MM_ADDR_RESET 32'h0

// DEBUG_S2MM_ADDR.ADDR - Indicates the Start Address
`define DMA_CSR_DEBUG_S2MM_ADDR_ADDR_WIDTH 32
`define DMA_CSR_DEBUG_S2MM_ADDR_ADDR_LSB 0
`define DMA_CSR_DEBUG_S2MM_ADDR_ADDR_MASK 32'hfc
`define DMA_CSR_DEBUG_S2MM_ADDR_ADDR_RESET 32'h0


`endif // __DMAREGS_VH