// Created with Corsair v1.0.2.dev0+894dec23
package DmaRegs_pkg;

parameter DMA_CSR_BASE_ADDR = 0;
parameter DMA_CSR_DATA_WIDTH = 32;
parameter DMA_CSR_ADDR_WIDTH = 8;

// DEBUG_CR
parameter DMA_CSR_DEBUG_CR_ADDR = 8'hf0;
parameter DMA_CSR_DEBUG_CR_RESET = 32'h0;

// DEBUG_CR.MM2S_LEN
parameter DMA_CSR_DEBUG_CR_MM2S_LEN_WIDTH = 8;
parameter DMA_CSR_DEBUG_CR_MM2S_LEN_LSB = 0;
parameter DMA_CSR_DEBUG_CR_MM2S_LEN_MASK = 32'hff;
parameter DMA_CSR_DEBUG_CR_MM2S_LEN_RESET = 8'h0;

// DEBUG_CR.MM2S_SIZE
parameter DMA_CSR_DEBUG_CR_MM2S_SIZE_WIDTH = 3;
parameter DMA_CSR_DEBUG_CR_MM2S_SIZE_LSB = 8;
parameter DMA_CSR_DEBUG_CR_MM2S_SIZE_MASK = 32'h700;
parameter DMA_CSR_DEBUG_CR_MM2S_SIZE_RESET = 3'h0;

// DEBUG_CR.MM2S_START
parameter DMA_CSR_DEBUG_CR_MM2S_START_WIDTH = 1;
parameter DMA_CSR_DEBUG_CR_MM2S_START_LSB = 12;
parameter DMA_CSR_DEBUG_CR_MM2S_START_MASK = 32'h1000;
parameter DMA_CSR_DEBUG_CR_MM2S_START_RESET = 1'h0;

// DEBUG_CR.S2MM_LEN
parameter DMA_CSR_DEBUG_CR_S2MM_LEN_WIDTH = 8;
parameter DMA_CSR_DEBUG_CR_S2MM_LEN_LSB = 16;
parameter DMA_CSR_DEBUG_CR_S2MM_LEN_MASK = 32'hff0000;
parameter DMA_CSR_DEBUG_CR_S2MM_LEN_RESET = 8'h0;

// DEBUG_CR.S2MM_SIZE
parameter DMA_CSR_DEBUG_CR_S2MM_SIZE_WIDTH = 3;
parameter DMA_CSR_DEBUG_CR_S2MM_SIZE_LSB = 24;
parameter DMA_CSR_DEBUG_CR_S2MM_SIZE_MASK = 32'h7000000;
parameter DMA_CSR_DEBUG_CR_S2MM_SIZE_RESET = 3'h0;

// DEBUG_CR.S2MM_START
parameter DMA_CSR_DEBUG_CR_S2MM_START_WIDTH = 1;
parameter DMA_CSR_DEBUG_CR_S2MM_START_LSB = 28;
parameter DMA_CSR_DEBUG_CR_S2MM_START_MASK = 32'h10000000;
parameter DMA_CSR_DEBUG_CR_S2MM_START_RESET = 1'h0;


// DEBUG_SR
parameter DMA_CSR_DEBUG_SR_ADDR = 8'hf4;
parameter DMA_CSR_DEBUG_SR_RESET = 32'h0;

// DEBUG_SR.MM2S_BUSY
parameter DMA_CSR_DEBUG_SR_MM2S_BUSY_WIDTH = 1;
parameter DMA_CSR_DEBUG_SR_MM2S_BUSY_LSB = 0;
parameter DMA_CSR_DEBUG_SR_MM2S_BUSY_MASK = 32'h1;
parameter DMA_CSR_DEBUG_SR_MM2S_BUSY_RESET = 1'h0;

// DEBUG_SR.S2MM_BUSY
parameter DMA_CSR_DEBUG_SR_S2MM_BUSY_WIDTH = 1;
parameter DMA_CSR_DEBUG_SR_S2MM_BUSY_LSB = 1;
parameter DMA_CSR_DEBUG_SR_S2MM_BUSY_MASK = 32'h2;
parameter DMA_CSR_DEBUG_SR_S2MM_BUSY_RESET = 1'h0;


// DEBUG_MM2S_ADDR
parameter DMA_CSR_DEBUG_MM2S_ADDR_ADDR = 8'hf8;
parameter DMA_CSR_DEBUG_MM2S_ADDR_RESET = 32'h0;

// DEBUG_MM2S_ADDR.ADDR
parameter DMA_CSR_DEBUG_MM2S_ADDR_ADDR_WIDTH = 32;
parameter DMA_CSR_DEBUG_MM2S_ADDR_ADDR_LSB = 0;
parameter DMA_CSR_DEBUG_MM2S_ADDR_ADDR_MASK = 32'hffffffff;
parameter DMA_CSR_DEBUG_MM2S_ADDR_ADDR_RESET = 32'h0;


// DEBUG_S2MM_ADDR
parameter DMA_CSR_DEBUG_S2MM_ADDR_ADDR = 8'hfc;
parameter DMA_CSR_DEBUG_S2MM_ADDR_RESET = 32'h0;

// DEBUG_S2MM_ADDR.ADDR
parameter DMA_CSR_DEBUG_S2MM_ADDR_ADDR_WIDTH = 32;
parameter DMA_CSR_DEBUG_S2MM_ADDR_ADDR_LSB = 0;
parameter DMA_CSR_DEBUG_S2MM_ADDR_ADDR_MASK = 32'hffffffff;
parameter DMA_CSR_DEBUG_S2MM_ADDR_ADDR_RESET = 32'h0;


endpackage