`ifndef _COEFFICIENT_SVH_
`define _COEFFICIENT_SVH_

package Coefficient;
    parameter real Alpha    = -1.586134342;
    parameter real Beta     = -0.052980118;
    parameter real Gama     =  0.882911076;
    parameter real Delta    =  0.443506852;
    parameter real K        = 1/(1.149604398);
endpackage

`endif // _COEFFICIENT_SVH_
