module Dwt97 #(
    parameter DataWidth = 16,
    parameter NumChannels = 1,
    parameter MaximumSideSize = 512
) (
    
);
    
endmodule