interface AxiStream (input clk);

endinterface //AxiStream